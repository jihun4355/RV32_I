// `timescale 1ns / 1ps
// module instr_mem (
//     input  logic [31:0] instr_rAddr,
//     output logic [31:0] instr_code
// );
//     logic [31:0] rom[0:63];

//     // initial begin
//     //     $readmemh("code2.txt", rom);
//     // end

//     initial begin
//         for (int i = 0; i < 64; i++) begin
//             rom[i] = 32'hffff_0000 + i;
//         end

// // // //////////////////////////////////////////////////////////////////////////////////////////
//         // // R-TYPE
//         // rom[0]  = 32'h004182B3;  //32'b0000_0000_0100_0001_1000_0010_1011_0011
//         // rom[1]  = 32'h409403B3;  //32'b0100_0000_1001_0100_0000_0011_1011_0011


// // // //////////////////////////////////////////////////////////////////////////////////////////

// //         // S-Type
// //         // 32'b imm(7bit) – rs2(5bit) – rs1(5bit) – funct3(3bit) – imm(5bit) - opcode(7bit)
// //         rom[2]  = 32'h00610223;  // sb x6, 7(x2) // 32'b0000000_00110_00010_010_00010_0100011; 
// //         rom[3]  = 32'h00811323;  // sh x8, 6(x2) // 32'b0000000_00000_00010_000_00111_0100011
// //         rom[4]  = 32'h00912323;  // sw x9, 6(x2) // 32'b0000000_01000_00010_001_01000_0100011
// //         rom[5]  = 32'h00610323;  // sb x6, 7(x2) // 32'b0000000_00011_00010_000_00010_0100011

// // //////////////////////////////////////////////////////////////////////////////////////////


//         // // IL-Type
//         // // // 32'b000000001100_00110_010_10101_0000011;
//         // rom[6]  = 32'h00C10083;  // lb x1, 12(x2) // 32'b 000000001100_00010_000_00001_0000011
//         // rom[7]  = 32'h00E11103;  // lh x2, 14(x2) // 32'b 000000001110_00010_001_00010_0000011
//         // rom[8]  = 32'h00C1_1283; // lw x5, 12(x2) // 32'b 000000001100_00010_010_00101_0000011
//         // rom[9]  = 32'h01214403;  // lbu x8, 18(x2) // 32'b 000000010010_00010_100_01000_0000011
//         // rom[10] = 32'h01414503;  // lhu x10, 20(x2) // 32'b 000000010100_00010_101_01010_0000011




//         // rom[1]  = 32'b000000001100_00010_000_00001_0000011;
//         // rom[2]  = 32'b000000001110_00010_001_00010_0000011;
//         // rom[3]  = 32'b000000001100_00010_010_00101_0000011;
//         // rom[4]  = 32'b000000010010_00010_100_01000_0000011;
//         // rom[5]  = 32'b000000010100_00010_101_01010_0000011;


//         // rom[0] = 32'h00C10083;  // lb  x1, 12(x2)
//         // rom[1] = 32'h00E11103;  // lh  x2, 14(x2)
//         // rom[2] = 32'h00C12283;  // lw  x5, 12(x2)
//         // rom[3] = 32'h01214403;  // lbu x8, 18(x2)
//         // rom[4] = 32'h01415503;  // lhu x10, 20(x2)



//         // rom[0] = 32'h00C10083;  // lb  x1, 12(x2)
//         // rom[1] = 32'h00E11103;  // lh  x2, 14(x2)
//         // rom[2] = 32'h00C11283;  // lw  x3, 12(x2)
//         // // rom[4] = 32'h00E12203;  // lbu x4, 14(x2)
//         // // rom[5] = 32'h00C12283;  // lhu x5, 12(x2)
//         // rom[3]  = 32'b000000010010_00010_100_01000_0000011;
//         // rom[4]  = 32'b000000010100_00010_101_01010_0000011;

// // rom[1] = 32'h00C10083;  // lb  x1, 12(x2)
// // rom[2] = 32'h00C11103;  // lh  x2, 12(x2)
// // rom[3] = 32'h00C11283;  // lw  x3, 12(x2)
// // rom[4] = 32'h00C12203;  // lbu x4, 12(x2)
// // rom[5] = 32'h00C12283;  // lhu x5, 12(x2)


// // // //         //////////////////////////////////////////////////////////////////////////////////////////


//         // // I_TYPE
//         // // 32'b000000001100_00110_000_01000_0010011;

//         // rom[0] = 32'h00A10113;  // addi x2, x2, 10  = (12)

//         // // 2. SLTI : x4 = (x2 < 10)? 1 : 0  
//         // rom[1] = 32'h00A12213;  // slti x4, x2, 10 = (0)
//         // // 000000001010_00010_010_00100_0010011

//         // // 3. SLTIU : x7 = (x2 < 14)? 1 : 0 (unsigned 비교)  = (1)
//         // rom[2] = 32'h00E13393;  // sltiu x7, x2, 14
//         // // 000000001110_00010_011_00111_0010011

//         // // 4. XORI : x8 = x2 ^ 5  = (9)
//         // rom[3] = 32'h00514413;  // xori x8, x2, 5

//         // // 5. ORI : x9 = x2 | 12  = (12)
//         // rom[4] = 32'h00C16493;  // ori x9, x2, 12
//         // // 000000001100_00010_110_01001_0010011

//         // // 6. ANDI : x10 = x2 & 7 = (4)
//         // rom[5] = 32'h00717513;  // andi x10, x2, 7
//         // // 000000000111_00010_111_01010_0010011

//         // // 7. SLLI : x13 = x2 << 2
//         // rom[6] = 32'h00211693;  // slli x13, x2, 2
//         // // 000000000010_00010_001_01101_0010011


//         // // 8. SRLI : x14 = x2 >> 1 (논리 시프트)
//         // rom[7] = 32'h00115713;  // srli x14, x2, 1
//         // // 000000000001_00010_101_01110_0010011

//         // // 9. SRAI : x15 = x2 >> 3 (산술 시프트)
//         // rom[8] = 32'h40315793;  // srai x15, x2, 3
//         // // 010000000011_00010_101_01111_0010011
        
// // //////////////////////////////////////////////////////////////////////////////////////////



// // // b-type
// //         // 32'b imm(7bit) – rs2(5bit) – rs1(5bit) – funct3(3bit) – imm(5bit) - opcode(7bit)
// //         // 1. BEQ: x1   == x1, 점프 (+8) -> rom[2]
// //         // Assembly: beq x1, x1, 12
        
// //         rom[1] = 32'b0000000_00001_00001_000_01100_1100011;

// //         // 2. BNE: x1 != x2, 점프 (+12) -> rom[4]
// //         // Assembly: bne x1, x2, 12
// //         rom[4] = 32'b0000000_00010_00001_001_01100_1100011;


// //         // 3. BLT: x1 < x2 (signed), 점프 (+16) -> rom[7]
// //         // Assembly: blt x1, x2, 12
// //         rom[7] = 32'b0000000_00010_00001_100_01100_1100011;



// //         // 4. BGE: x2 >= x1 (signed), 점프 (+20) -> rom[12]
// //         // Assembly: bge x2, x1, 12
// //         rom[10] = 32'b0000000_00001_00010_101_01100_1100011;



// //         // 5. BLTU: x3 < x4 (unsigned), 점프 (+24) -> rom[18]
// //         // Assembly: bltu x3, x4, 12
// //         rom[13] = 32'b0000000_00100_00011_110_01100_1100011; 



// //         // 6. BGEU: x4 >= x3 (unsigned), 점프 (+28) -> rom[25]
// //         // Assembly: bgeu x4, x3, 12

// //         rom[16] = 32'b0000000_00011_00100_111_01100_1100011; 
        

//         // rom[1]  = 32'h00208663; // beq  x1, x1, 12
//         // rom[4]  = 32'h00209663; // bne  x1, x2, 12
//         // rom[7]  = 32'h0020C663; // blt  x1, x2, 12
//         // rom[10] = 32'h00115663; // bge  x2, x1, 12
//         // rom[13] = 32'h0041E663; // bltu x3, x4, 12
//         // rom[16] = 32'h00327663; // bgeu x4, x3, 12


// // //////////////////////////////////////////////////////////////////////////////////////////

//     //    // U_TYPE

        
//     //     rom[4] = 32'b00010000000000000000_00100_0110111; // lui x4, 0x10000 // rom[4] = 32'h00010437; // lui   x4, 0x10000
//     //     rom[5] = 32'b00010000000000000000_00101_0010111; // auipc x5, 0x10000 // rom[5] = 32'h00010517; // auipc x5, 0x10000

        
        

// // //////////////////////////////////////////////////////////////////////////////////////////


//         // J-  type
//             rom [0]  = 32'b0000000000100_00010_000_01000_1100111; // JALR // rom[0] = 32'h00410067; // jalr x8, x2, 4
//             rom [4]  = 32'b00000000000000000100_00100_1101111;    // JAL  // rom[4] = 32'h0040026F; // jal  x4, 4

//     //    //////////////////////////////////////////////////////////////////////////////////////////

            
//     //     //R-TYPE
//     //     rom[0]  = 32'h004182B3;  // add  x5, x3, x4
//     //     rom[1]  = 32'h409403B3;  // sub  x7, x8, x9

//     //     //////////////////////////////////////////////////////////////////////////////////////////
//     //     // S-TYPE
//     //     rom[2]  = 32'h00610223;  // sb x6, 7(x2)
//     //     rom[3]  = 32'h00811323;  // sh x8, 6(x2)
//     //     rom[4]  = 32'h00912323;  // sw x9, 6(x2)
//     //     rom[5]  = 32'h00610323;  // sb x6, 7(x2)

//     //     //////////////////////////////////////////////////////////////////////////////////////////
//     //     // IL-TYPE (LOAD)
//     //     rom[6]  = 32'h00C10083;  // lb  x1, 12(x2)
//     //     rom[7]  = 32'h00E11103;  // lh  x2, 14(x2)
//     //     rom[8]  = 32'h00C11283;  // lw  x5, 12(x2)
//     //     rom[9]  = 32'h01214403;  // lbu x8, 18(x2)
//     //     rom[10] = 32'h01414503;  // lhu x10, 20(x2)

//     //     //////////////////////////////////////////////////////////////////////////////////////////
//     //     // I-TYPE
//     //     rom[12] = 32'h00A10113;  // addi  x2, x2, 10
//     //     rom[13] = 32'h00A12213;  // slti  x4, x2, 10
//     //     rom[14] = 32'h00E13393;  // sltiu x7, x2, 14
//     //     rom[15] = 32'h00514413;  // xori  x8, x2, 5
//     //     rom[16] = 32'h00C16493;  // ori   x9, x2, 12
//     //     rom[17] = 32'h00717513;  // andi  x10, x2, 7
//     //     rom[18] = 32'h00211693;  // slli  x13, x2, 2
//     //     rom[19] = 32'h00115713;  // srli  x14, x2, 1
//     //     rom[20] = 32'h40315793;  // srai  x15, x2, 3

//     //     //////////////////////////////////////////////////////////////////////////////////////////

//     //     // B-TYPE (branch offset = 12)
//     //     rom[21] = 32'h00208663;   // beq  x1, x1, 12
//     //     rom[22] = 32'h00209663; // bne  x1, x2, 12
//     //     rom[23] = 32'h0020C663;   // blt  x1, x2, 12
//     //     rom[24] = 32'h00115663;  // bge  x2, x1, 12
//     //     rom[25] = 32'h0041E663;  // bltu x3, x4, 12
//     //     rom[26] = 32'h00327663;  // bgeu x4, x3, 12



//     // //     // //////////////////////////////////////////////////////////////////////////////////////////



// // 2진수(4bit)	16진수
// // 0000	0
// // 0001	1
// // 0010	2
// // 0011	3
// // 0100	4
// // 0101	5
// // 0110	6
// // 0111	7
// // 1000	8
// // 1001	9
// // 1010	A
// // 1011	B
// // 1100	C
// // 1101	D
// // 1110	E
// // 1111	F


// //    // x4 → 00100
// //
// //    // x8 → 01000
// //
// //    // x12 → 01100
// //
// //    // x16 → 10000                           
//     end

//     assign instr_code = rom[instr_rAddr[31:2]];

// endmodule







































`timescale 1ns / 1ps

module instr_mem (
    input  logic [31:0] instr_rAddr,
    output logic [31:0] instr_code
);
    logic [31:0] rom[0:200];

    initial begin
        $readmemh("code_0929_exam0.mem", rom);


        // // R-TYPE
        // rom[0] = 32'b0000_0000_0100_0001_1000_0010_1011_0011;
        // rom[1] = 32'b0100_0000_1001_0100_0000_0011_1011_0011;
        // rom[2] = 32'b0000_0000_0111_0100_1111_0000_1011_0011;
        // rom[3] = 32'b0000_0000_0001_0100_1000_0100_1011_0011;
        // rom[4] = 32'b0000_0000_0010_0010_0100_0011_1011_0011;
        // rom[5] = 32'b0000_0000_0110_0011_1001_0010_1011_0011;
        // rom[6] = 32'b0000_0000_1000_0010_1100_0100_1011_0011;
        // rom[7] = 32'b0100_0000_1001_0001_1001_0001_1011_0011;
        // rom[8] = 32'b0000_0000_0100_0100_1011_0001_1011_0011;
        // rom[9] = 32'b0000_0000_0011_0011_0100_0100_1011_0011;

        // add 2 + 3 = 5
        // sub 3 - 4 = -1
        // sll 4 << 5 = 128
        // srl 5 >> 6 = 0
        // sra 6 >>> 7 = 0
        // slt 7 < 8  = 1
        // sltu 8 < 9 = 1
        // xor 9 ^ 10 = 3
        // or 10 | 11 = 11
        // and 11 & 12 = 8

        // rom[0] = 32'h003100b3;
        // rom[1] = 32'h40418133;
        // rom[2] = 32'h005211b3;
        // rom[3] = 32'h0062d233;
        // rom[4] = 32'h407352b3;
        // rom[5] = 32'h0083a333;
        // rom[6] = 32'h009433b3;
        // rom[7] = 32'h00a4c433;
        // rom[8] = 32'h00b564b3;
        // rom[9] = 32'h00c5f533;



        // ADD    4, 3, 5    0000_0000_0100_0001_1000_0010_1011_0011 4 + 3 = 7
        // SUB    9, 8, 7    0100_0000_1001_0100_0000_0011_1011_0011 8 - 9 = -1
        // AND    7, 9, 1    0000_0000_0111_0100_1111_0000_1011_0011 9 & 7 = 1
        // OR     1, 8, 9    0000_0000_0001_0100_1000_0100_1011_0011 1 | 8 = 9
        // SLT    2, 4, 6    0000_0000_0010_0010_0100_0011_1011_0011 x4 < x6 ? 1 : 0 = 0
        // SLL    6, 7, 5    0000_0000_0110_0011_1001_0010_1011_0011
        // SRL    8, 5, 4    0000_0000_1000_0010_1100_0100_1011_0011
        // SRA    9, 3, 2    0100_0000_1001_0001_1001_0001_1011_0011
        // SLT(U) 4, 9, 3    0000_0000_0100_0100_1011_0001_1011_0011
        // XOR    3, 6, 8    0000_0000_0011_0011_0100_0100_1011_0011


        // // S-Type
        // rom[3]  = 32'h00811323;  // sh x8, 6(x2)
        // rom[4]  = 32'h00912323;  // sw x9, 6(x2)
        // rom[5]  = 32'h00610323;  // sb x6, 6(x2)

        // // IL-Type
        // rom[1] = 32'h00130083;  // lb x1, 1(x6)
        // rom[2] = 32'h00231103;  // lh x2, 2(x6)
        // rom[3] = 32'h00332183;  // lw x3, 3(x6)
        // rom[4] = 32'h00434203;  // lbu x4, 4(x6)
        // rom[5] = 32'h0053d283;  // lhu x5, 5(x6)


        // // I_TYPE
        // // 1. ADDI : x2 = x2 + 10
        // rom[0] = 32'h00A10113;  // addi x2, x2, 10  = (12)

        // // 2. SLTI : x4 = (x2 < 10)? 1 : 0  
        // rom[1] = 32'h00A12213;  // slti x4, x2, 10 = (0)

        // // 3. SLTIU : x7 = (x2 < 14)? 1 : 0 (unsigned 비교)  = (1)
        // rom[2] = 32'h00E13393;  // sltiu x7, x2, 14

        // // 4. XORI : x8 = x2 ^ 5  = (9)
        // rom[3] = 32'h00514413;  // xori x8, x2, 5

        // // 5. ORI : x9 = x2 | 12  = (12)
        // rom[4] = 32'h00C16493;  // ori x9, x2, 12

        // // 6. ANDI : x10 = x2 & 7 = (4)
        // rom[5] = 32'h00717513;  // andi x10, x2, 7

        // // 7. SLLI : x13 = x2 << 2
        // rom[6] = 32'h00211693;  // slli x13, x2, 2

        // // 8. SRLI : x14 = x2 >> 1 (논리 시프트)
        // rom[7] = 32'h00115713;  // srli x14, x2, 1
 
        // // 9. SRAI : x15 = x2 >> 3 (산술 시프트)
        // rom[8] = 32'h40315793;  // srai x15, x2, 3



        // B-TYPE

        // rom[0] = 32'h00210463;    // BEQ  x2, x2, 8    if(rs1 == rs2) PC += imm
        // rom[1] = 32'b0000_0000_0100_0001_1000_0010_1011_0011; // add
        // rom[2] = 32'h001114631;   // BNE  x1, x2, 8   if(rs1 != rs2) PC += imm
        // rom[3] = 32'b0000_0000_0100_0001_1000_0010_1011_0011; // add
        // rom[4] = 32'h0020c463;   // BLT  x2, x1, 8   if(rs1 < rs2) PC += imm
        // rom[5] = 32'b0000_0000_0100_0001_1000_0010_1011_0011; // add
        // rom[6] = 32'h0023d463;   // BGE  x2, x7, 8   if(rs1 >= rs2) PC += imm  
        // rom[7] = 32'b0000_0000_0100_0001_1000_0010_1011_0011; // add
        // rom[8] = 32'h00416463;   // BLTU x4, x2, 8    if(rs1 < rs2) PC += imm
        // rom[9] = 32'b0000_0000_0100_0001_1000_0010_1011_0011; // add
        // rom[10] = 32'h00547463;   // BGEU x5, x8, 8   if(rs1 >= rs2) PC += imm


        // // U_TYPE
        // rom[0] = 32'b0000_0000_0000_0000_0010_00001_0110111;  // LUI  x1 = 2  rd = imm
        // rom[1] = 32'b0000_0000_0000_0000_0100_00100_0010111;  // AUIPC  x3 = 4 + 4 = 8 rd = PC + imm

        // J_TYPE
        rom[0] = 32'h0061_02E7;  // JARL x5, x2, 6 
        // rom[1] = 32'h0080_02EF;  // JAL  x5, 8
        rom[2] = 32'h0080_02EF;  // JAL  x5, 8

    end

    assign instr_code = rom[instr_rAddr[31:2]];

endmodule

























